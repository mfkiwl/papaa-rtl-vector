module vv_fsm
  # (parameter N=4)
    (input clk,
     input rst,
     input start,
     output reg [$clog2(N)-1:0] rd_addr,
     output reg mem_wr_en,
     output reg [$clog2(N)-1:0] wr_addr,
     output reg init
     );


// insert code here

endmodule
